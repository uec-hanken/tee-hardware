module inv_mixw (
	input	[31:0]	w,
	output	[31:0]	out
);

assign out[31] = w[30]^w[29]^w[28]^w[23]^w[22]^w[20]^w[15]^w[13]^w[12]^w[7] ^w[4];
assign out[30] = w[31]^w[29]^w[28]^w[27]^w[23]^w[22]^w[21]^w[19]^w[15]^w[14]^w[12]^w[11]^w[7] ^w[6] ^w[3];
assign out[29] = w[30]^w[28]^w[27]^w[26]^w[23]^w[22]^w[21]^w[20]^w[18]^w[14]^w[13]^w[11]^w[10]^w[7] ^w[6]^w[5]^w[2];
assign out[28] = w[29]^w[27]^w[26]^w[25]^w[23]^w[22]^w[21]^w[20]^w[19]^w[17]^w[15]^w[13]^w[12]^w[10]^w[9]^w[6]^w[5]^w[4]^w[1];
assign out[27] = w[30]^w[29]^w[26]^w[25]^w[24]^w[21]^w[19]^w[18]^w[16]^w[15]^w[14]^w[13]^w[11]^w[9] ^w[8]^w[7]^w[5]^w[3]^w[0];
assign out[26] = w[30]^w[25]^w[24]^w[23]^w[22]^w[18]^w[17]^w[14]^w[10]^w[8] ^w[7] ^w[6] ^w[2];
assign out[25] = w[29]^w[24]^w[23]^w[22]^w[21]^w[17]^w[16]^w[15]^w[13]^w[9] ^w[6] ^w[5] ^w[1];
assign out[24] = w[31]^w[30]^w[29]^w[23]^w[21]^w[16]^w[14]^w[13]^w[8] ^w[5] ^w[0];
assign out[23] = w[31]^w[28]^w[22]^w[21]^w[20]^w[15]^w[14]^w[12]^w[7] ^w[5] ^w[4];
assign out[22] = w[31]^w[30]^w[27]^w[23]^w[21]^w[20]^w[19]^w[15]^w[14]^w[13]^w[11]^w[7] ^w[6] ^w[4]^w[3];
assign out[21] = w[31]^w[30]^w[29]^w[26]^w[22]^w[20]^w[19]^w[18]^w[15]^w[14]^w[13]^w[12]^w[10]^w[6]^w[5]^w[3]^w[2];
assign out[20] = w[30]^w[29]^w[28]^w[25]^w[21]^w[19]^w[18]^w[17]^w[15]^w[14]^w[13]^w[12]^w[11]^w[9]^w[7]^w[5]^w[4]^w[2]^w[1];
assign out[19] = w[31]^w[29]^w[27]^w[24]^w[22]^w[21]^w[18]^w[17]^w[16]^w[13]^w[11]^w[10]^w[8] ^w[7]^w[6]^w[5]^w[3]^w[1]^w[0];
assign out[18] = w[31]^w[30]^w[26]^w[22]^w[17]^w[16]^w[15]^w[14]^w[10]^w[9] ^w[6] ^w[2] ^w[0];
assign out[17] = w[30]^w[29]^w[25]^w[21]^w[16]^w[15]^w[14]^w[13]^w[9] ^w[8] ^w[7] ^w[5] ^w[1];
assign out[16] = w[29]^w[24]^w[23]^w[22]^w[21]^w[15]^w[13]^w[8] ^w[6] ^w[5] ^w[0];
assign out[15] = w[31]^w[29]^w[28]^w[23]^w[20]^w[14]^w[13]^w[12]^w[7] ^w[6] ^w[4];
assign out[14] = w[31]^w[30]^w[28]^w[27]^w[23]^w[22]^w[19]^w[15]^w[13]^w[12]^w[11]^w[7] ^w[6] ^w[5]^w[3];
assign out[13] = w[30]^w[29]^w[27]^w[26]^w[23]^w[22]^w[21]^w[18]^w[14]^w[12]^w[11]^w[10]^w[7] ^w[6]^w[5]^w[4]^w[2];
assign out[12] = w[31]^w[29]^w[28]^w[26]^w[25]^w[22]^w[21]^w[20]^w[17]^w[13]^w[11]^w[10]^w[9] ^w[7]^w[6]^w[5]^w[4]^w[3]^w[1];
assign out[11] = w[31]^w[30]^w[29]^w[27]^w[25]^w[24]^w[23]^w[21]^w[19]^w[16]^w[14]^w[13]^w[10]^w[9]^w[8]^w[5]^w[3]^w[2]^w[0];
assign out[10] = w[30]^w[26]^w[24]^w[23]^w[22]^w[18]^w[14]^w[9] ^w[8] ^w[7] ^w[6] ^w[2] ^w[1];
assign out[9]  = w[31]^w[29]^w[25]^w[22]^w[21]^w[17]^w[13]^w[8] ^w[7] ^w[6] ^w[5] ^w[1] ^w[0];
assign out[8]  = w[30]^w[29]^w[24]^w[21]^w[16]^w[15]^w[14]^w[13]^w[7] ^w[5] ^w[0];
assign out[7]  = w[31]^w[30]^w[28]^w[23]^w[21]^w[20]^w[15]^w[12]^w[6] ^w[5] ^w[4];
assign out[6]  = w[31]^w[30]^w[29]^w[27]^w[23]^w[22]^w[20]^w[19]^w[15]^w[14]^w[11]^w[7] ^w[5] ^w[4] ^w[3];
assign out[5]  = w[31]^w[30]^w[29]^w[28]^w[26]^w[22]^w[21]^w[19]^w[18]^w[15]^w[14]^w[13]^w[10]^w[6] ^w[4]^w[3]^w[2];
assign out[4]  = w[31]^w[30]^w[29]^w[28]^w[27]^w[25]^w[23]^w[21]^w[20]^w[18]^w[17]^w[14]^w[13]^w[12]^w[9]^w[5]^w[3]^w[2]^w[1];
assign out[3]  = w[29]^w[27]^w[26]^w[24]^w[23]^w[22]^w[21]^w[19]^w[17]^w[16]^w[15]^w[13]^w[11]^w[8] ^w[6]^w[5]^w[2]^w[1]^w[0];
assign out[2]  = w[31]^w[30]^w[26]^w[25]^w[22]^w[18]^w[16]^w[15]^w[14]^w[10]^w[6] ^w[1] ^w[0];
assign out[1]  = w[31]^w[30]^w[29]^w[25]^w[24]^w[23]^w[21]^w[17]^w[14]^w[13]^w[9] ^w[5] ^w[0];
assign out[0]  = w[31]^w[29]^w[24]^w[22]^w[21]^w[16]^w[13]^w[8] ^w[7] ^w[6] ^w[5];

endmodule

module inv_mixcolumns (
	input	[127:0]	data,
	output	[127:0]	out
);

inv_mixw u3 (
	.w		(data[127:96]),
	.out	(out[127:96])
);

inv_mixw u2 (
	.w		(data[95:64]),
	.out	(out[95:64])
);

inv_mixw u1 (
	.w		(data[63:32]),
	.out	(out[63:32])
);

inv_mixw u0 (
	.w		(data[31:0]),
	.out	(out[31:0])
);

endmodule
